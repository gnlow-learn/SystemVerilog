module helloworld;
    initial begin
        $display("Hello, World!");
    end
endmodule
